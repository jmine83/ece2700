`timescale 1ns / 1ps

module Multiplier_T();

	reg S7_s, S6_s, S5_s, S4_s, S3_s, S2_s, S1_s, S0_s;
	wire [7:0] PR_s;

	Multiplier test(S7_s, S6_s, S5_s, S4_s, S3_s, S2_s, S1_s, S0_s, PR_s);

	initial begin
		S7_s <= 0; S6_s <= 0; S5_s <= 0; S4_s <= 0; S3_s <= 0; S2_s <= 0; S1_s <= 0; S0_s <= 0; // 0 * 0 = 0
		#10 S7_s <= 0; S6_s <= 0; S5_s <= 1; S4_s <= 0;  S3_s <= 0; S2_s <= 0; S1_s <= 1; S0_s <= 1; // 2 * 3 = 6
		#10 S7_s <= 0; S6_s <= 0; S5_s <= 1; S4_s <= 1;  S3_s <= 0; S2_s <= 0; S1_s <= 1; S0_s <= 1; // 3 * 3 = 9
		#10 S7_s <= 0; S6_s <= 1; S5_s <= 0; S4_s <= 1;  S3_s <= 0; S2_s <= 0; S1_s <= 1; S0_s <= 0; // 5 * 2 = 10
		#10 S7_s <= 1; S6_s <= 0; S5_s <= 0; S4_s <= 0;  S3_s <= 0; S2_s <= 1; S1_s <= 0; S0_s <= 0; // 8 * 4 = 32
		#10 S7_s <= 1; S6_s <= 0; S5_s <= 0; S4_s <= 1;  S3_s <= 0; S2_s <= 1; S1_s <= 1; S0_s <= 0; // 9 * 6 = 54
		#10 S7_s <= 1; S6_s <= 0; S5_s <= 1; S4_s <= 1;  S3_s <= 1; S2_s <= 0; S1_s <= 0; S0_s <= 1; // 11 * 9 = 99
		#10 S7_s <= 1; S6_s <= 0; S5_s <= 1; S4_s <= 0;  S3_s <= 1; S2_s <= 0; S1_s <= 1; S0_s <= 0; // 10 * 10 = 100
		#10 S7_s <= 1; S6_s <= 1; S5_s <= 0; S4_s <= 1;  S3_s <= 1; S2_s <= 0; S1_s <= 0; S0_s <= 0; // 13 * 8 = 104
		#10 S7_s <= 1; S6_s <= 1; S5_s <= 0; S4_s <= 0;  S3_s <= 1; S2_s <= 0; S1_s <= 1; S0_s <= 0; // 12 * 10 = 120
		#10 S7_s <= 1; S6_s <= 1; S5_s <= 0; S4_s <= 0;  S3_s <= 1; S2_s <= 1; S1_s <= 0; S0_s <= 0; // 12 * 12 = 144
		#10 S7_s <= 1; S6_s <= 1; S5_s <= 1; S4_s <= 1;  S3_s <= 1; S2_s <= 0; S1_s <= 1; S0_s <= 1; // 15 * 11 = 165
		#10 S7_s <= 1; S6_s <= 1; S5_s <= 1; S4_s <= 1;  S3_s <= 1; S2_s <= 1; S1_s <= 1; S0_s <= 0; // 15 * 14 = 210
		#10 S7_s <= 1; S6_s <= 1; S5_s <= 1; S4_s <= 1;  S3_s <= 1; S2_s <= 1; S1_s <= 1; S0_s <= 1; // 15 * 15 = 225
	end
	
endmodule
